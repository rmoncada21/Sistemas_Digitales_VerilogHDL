module FFD_reset_sync(
    
);

endmodule