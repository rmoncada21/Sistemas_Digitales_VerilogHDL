// Circuito del ejercicio 4.1 modelado por comportamiento
// Modelado por comportamiento
module circuito_mpc (A, B, C, D, F1, F2);
    input A, B, C, D;
    output F1, F2;

endmodule