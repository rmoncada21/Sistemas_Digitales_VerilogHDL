module reg4_paralell_load_with_FFD;
    // puertos del test

    // variables del test

    // instanciación del uut/dut

    // task del testbench

    // inicialización de las variables
endmodule