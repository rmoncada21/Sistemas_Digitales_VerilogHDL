// Modelado por flujo de datos

module circuito_mfd(A, B, C, D, F1, F2);
    input A, B, C, D;
    output F1, F2;
    
endmodule