`timescale 1ns/1ps 
module g_and(input A, input B, output Y);
    assign Y = A & B;  // Operación AND
endmodule
